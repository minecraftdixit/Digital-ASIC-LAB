`timescale 1ns / 1ps
 
module Adder (
  input [15:0] in1,
  input [15:0] in2,
  output [15:0] sum
);

assign sum = in1 + in2;

endmodule : Adder
